`include "design.sv"
`include "multiplier_trans.sv"
`include "multiplier_gen.sv"
`include "multiplier_intf.sv"
`include "multiplier_bfm.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "multiplier_cov.sv"
`include "multiplier_env.sv"
`include "multiplier_test.sv"
`include "tb_multiplier_top_tb.sv"



